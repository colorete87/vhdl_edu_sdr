-- libraries
library ieee;
use ieee.std_logic_1164.all;

entity top_uart is
end entity top_uart;


architecture rtl of top_uart is
begin
end architecture;
